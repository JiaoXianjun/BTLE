// Author: Xianjun Jiao <putaoshu@msn.com>
// SPDX-FileCopyrightText: 2024 Xianjun Jiao
// SPDX-License-Identifier: Apache-2.0 license

// To generate test vector:
// Create bit_repeat_upsample_test_input.txt with 1 bit (0 or 1) per line
// Run verilog simulation:
// iverilog -o bit_repeat_upsample_tb bit_repeat_upsample_tb.v bit_repeat_upsample.v
// vvp bit_repeat_upsample_tb
// Then remove the "// address " comment lines form file generated by writememh()
// grep -v // bit_repeat_upsample_test_output.txt > new.txt
// Each bit in the _test_input.txt will be repeated 8 times

// ATTENTION: NUM_BIT_INPUT needs to be equal to the number of lines in bit_repeat_upsample_test_input.txt
`timescale 1ns / 1ps
module bit_repeat_upsample_tb #
(
  parameter SAMPLE_PER_SYMBOL = 8,
  parameter NUM_BIT_INPUT = 11
) (
);

reg clk;
reg rst;

reg [0:0] bit_repeat_upsample_test_input_mem [0:4095];
reg [0:0] bit_repeat_upsample_test_output_mem [0:4095];
initial begin
  $dumpfile("bit_repeat_upsample_tb.vcd");
  $dumpvars;
  $readmemh("bit_repeat_upsample_test_input.txt", bit_repeat_upsample_test_input_mem);

  clk = 0;
  rst = 0;
  
  #200 rst = 1;

  #200 rst = 0;
end

always begin
  #((1000.0/16.0)/2.0) clk = !clk; //16MHz
end

reg bit;
reg bit_valid;
reg bit_valid_last;

wire bit_upsample;
wire bit_upsample_valid;
wire bit_upsample_valid_last;

// test process
reg [31:0] clk_count;
reg [31:0] info_bit_count;
reg [31:0] bit_out_count;
always @ (posedge clk) begin
  if (rst) begin
    bit <= 0;
    bit_valid <= 0;

    clk_count <= 1;
    info_bit_count <= 0;
    bit_out_count <= 0;
  end else begin
    clk_count <= clk_count + 1;

    if (clk_count[3:0] == 0) begin // speed 1M
      if (info_bit_count < NUM_BIT_INPUT) begin
        bit <= bit_repeat_upsample_test_input_mem[info_bit_count];
        bit_valid <= 1;
        // $display("%h", bit_repeat_upsample_test_input_mem[info_bit_count]);
        if (info_bit_count == (NUM_BIT_INPUT-1)) begin
          bit_valid_last <= 1;
        end
      end
      info_bit_count <= info_bit_count + 1;
    end else begin
      bit_valid <= 0;
      bit_valid_last <= 0;
    end

    if (info_bit_count == (NUM_BIT_INPUT+30)) begin
      $display("%d input", NUM_BIT_INPUT);
      $display("%d output", bit_out_count);
      $writememh("bit_repeat_upsample_test_output.txt", bit_repeat_upsample_test_output_mem, 0, bit_out_count-1);
      $display("Please compare bit_repeat_upsample_test_output.txt and bit_repeat_upsample_test_input.txt");
      $finish;
    end

    // record the result
    if (bit_upsample_valid) begin
      bit_repeat_upsample_test_output_mem[bit_out_count] <= bit_upsample;
      bit_out_count <= bit_out_count + 1;
    end
  end
end

bit_repeat_upsample # (
  .SAMPLE_PER_SYMBOL(SAMPLE_PER_SYMBOL)        
) bit_repeat_upsample_i (
  .clk(clk),
  .rst(rst),

  .phy_bit(bit),
  .bit_valid(bit_valid),
  .bit_valid_last(bit_valid_last),

  .bit_upsample(bit_upsample),
  .bit_upsample_valid(bit_upsample_valid),
  .bit_upsample_valid_last(bit_upsample_valid_last)
);

endmodule

